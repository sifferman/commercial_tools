module tb;
    initial begin
        $display("Hello, World!");
        $finish;
    end
endmodule
